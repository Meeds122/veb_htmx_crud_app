module main

import veb
import time

fn main() {
	println('Hello World!')
}
